//TESTED
module Mux_Weight(In, Select, Out);

parameter OUT_SIZE = 133;
parameter SEL_SIZE = 112;
parameter SEL_BIT  = 7;

input       [OUT_SIZE*SEL_SIZE-1:0]     In;
input       [SEL_BIT-1:0]               Select;
output  reg [OUT_SIZE-1:0]              Out;

always@(Select) begin
    case(Select)
        default:    Out = In[OUT_SIZE*1-1:OUT_SIZE*0];
        7'd1:       Out = In[OUT_SIZE*2-1:OUT_SIZE*1];
        7'd2:       Out = In[OUT_SIZE*3-1:OUT_SIZE*2];
        7'd3:       Out = In[OUT_SIZE*4-1:OUT_SIZE*3];
        7'd4:       Out = In[OUT_SIZE*5-1:OUT_SIZE*4];
        7'd5:       Out = In[OUT_SIZE*6-1:OUT_SIZE*5];
        7'd6:       Out = In[OUT_SIZE*7-1:OUT_SIZE*6];
        7'd7:       Out = In[OUT_SIZE*8-1:OUT_SIZE*7];
        7'd8:       Out = In[OUT_SIZE*9-1:OUT_SIZE*8];
        7'd9:       Out = In[OUT_SIZE*10-1:OUT_SIZE*9];
        7'd10:      Out = In[OUT_SIZE*11-1:OUT_SIZE*10];
        7'd11:      Out = In[OUT_SIZE*12-1:OUT_SIZE*11];
        7'd12:      Out = In[OUT_SIZE*13-1:OUT_SIZE*12];
        7'd13:      Out = In[OUT_SIZE*14-1:OUT_SIZE*13];
        7'd14:      Out = In[OUT_SIZE*15-1:OUT_SIZE*14];
        7'd15:      Out = In[OUT_SIZE*16-1:OUT_SIZE*15];
        7'd16:      Out = In[OUT_SIZE*17-1:OUT_SIZE*16];
        7'd17:      Out = In[OUT_SIZE*18-1:OUT_SIZE*17];
        7'd18:      Out = In[OUT_SIZE*19-1:OUT_SIZE*18];
        7'd19:      Out = In[OUT_SIZE*20-1:OUT_SIZE*19];
        7'd20:      Out = In[OUT_SIZE*21-1:OUT_SIZE*20];
        7'd21:      Out = In[OUT_SIZE*22-1:OUT_SIZE*21];
        7'd22:      Out = In[OUT_SIZE*23-1:OUT_SIZE*22];
        7'd23:      Out = In[OUT_SIZE*24-1:OUT_SIZE*23];
        7'd24:      Out = In[OUT_SIZE*25-1:OUT_SIZE*24];
        7'd25:      Out = In[OUT_SIZE*26-1:OUT_SIZE*25];
        7'd26:      Out = In[OUT_SIZE*27-1:OUT_SIZE*26];
        7'd27:      Out = In[OUT_SIZE*28-1:OUT_SIZE*27];
        7'd28:      Out = In[OUT_SIZE*29-1:OUT_SIZE*28];
        7'd29:      Out = In[OUT_SIZE*30-1:OUT_SIZE*29];
        7'd30:      Out = In[OUT_SIZE*31-1:OUT_SIZE*30];
        7'd31:      Out = In[OUT_SIZE*32-1:OUT_SIZE*31];
        7'd32:      Out = In[OUT_SIZE*33-1:OUT_SIZE*32];
        7'd33:      Out = In[OUT_SIZE*34-1:OUT_SIZE*33];
        7'd34:      Out = In[OUT_SIZE*35-1:OUT_SIZE*34];
        7'd35:      Out = In[OUT_SIZE*36-1:OUT_SIZE*35];
        7'd36:      Out = In[OUT_SIZE*37-1:OUT_SIZE*36];
        7'd37:      Out = In[OUT_SIZE*38-1:OUT_SIZE*37];
        7'd38:      Out = In[OUT_SIZE*39-1:OUT_SIZE*38];
        7'd39:      Out = In[OUT_SIZE*40-1:OUT_SIZE*39];
        7'd40:      Out = In[OUT_SIZE*41-1:OUT_SIZE*40];
        7'd41:      Out = In[OUT_SIZE*42-1:OUT_SIZE*41];
        7'd42:      Out = In[OUT_SIZE*43-1:OUT_SIZE*42];
        7'd43:      Out = In[OUT_SIZE*44-1:OUT_SIZE*43];
        7'd44:      Out = In[OUT_SIZE*45-1:OUT_SIZE*44];
        7'd45:      Out = In[OUT_SIZE*46-1:OUT_SIZE*45];
        7'd46:      Out = In[OUT_SIZE*47-1:OUT_SIZE*46];
        7'd47:      Out = In[OUT_SIZE*48-1:OUT_SIZE*47];
        7'd48:      Out = In[OUT_SIZE*49-1:OUT_SIZE*48];
        7'd49:      Out = In[OUT_SIZE*50-1:OUT_SIZE*49];
        7'd50:      Out = In[OUT_SIZE*51-1:OUT_SIZE*50];
        7'd51:      Out = In[OUT_SIZE*52-1:OUT_SIZE*51];
        7'd52:      Out = In[OUT_SIZE*53-1:OUT_SIZE*52];
        7'd53:      Out = In[OUT_SIZE*54-1:OUT_SIZE*53];
        7'd54:      Out = In[OUT_SIZE*55-1:OUT_SIZE*54];
        7'd55:      Out = In[OUT_SIZE*56-1:OUT_SIZE*55];
        7'd56:      Out = In[OUT_SIZE*57-1:OUT_SIZE*56];
        7'd57:      Out = In[OUT_SIZE*58-1:OUT_SIZE*57];
        7'd58:      Out = In[OUT_SIZE*59-1:OUT_SIZE*58];
        7'd59:      Out = In[OUT_SIZE*60-1:OUT_SIZE*59];
        7'd60:      Out = In[OUT_SIZE*61-1:OUT_SIZE*60];
        7'd61:      Out = In[OUT_SIZE*62-1:OUT_SIZE*61];
        7'd62:      Out = In[OUT_SIZE*63-1:OUT_SIZE*62];
        7'd63:      Out = In[OUT_SIZE*64-1:OUT_SIZE*63];
        7'd64:      Out = In[OUT_SIZE*65-1:OUT_SIZE*64];
        7'd65:      Out = In[OUT_SIZE*66-1:OUT_SIZE*65];
        7'd66:      Out = In[OUT_SIZE*67-1:OUT_SIZE*66];
        7'd67:      Out = In[OUT_SIZE*68-1:OUT_SIZE*67];
        7'd68:      Out = In[OUT_SIZE*69-1:OUT_SIZE*68];
        7'd69:      Out = In[OUT_SIZE*70-1:OUT_SIZE*69];
        7'd70:      Out = In[OUT_SIZE*71-1:OUT_SIZE*70];
        7'd71:      Out = In[OUT_SIZE*72-1:OUT_SIZE*71];
        7'd72:      Out = In[OUT_SIZE*73-1:OUT_SIZE*72];
        7'd73:      Out = In[OUT_SIZE*74-1:OUT_SIZE*73];
        7'd74:      Out = In[OUT_SIZE*75-1:OUT_SIZE*74];
        7'd75:      Out = In[OUT_SIZE*76-1:OUT_SIZE*75];
        7'd76:      Out = In[OUT_SIZE*77-1:OUT_SIZE*76];
        7'd77:      Out = In[OUT_SIZE*78-1:OUT_SIZE*77];
        7'd78:      Out = In[OUT_SIZE*79-1:OUT_SIZE*78];
        7'd79:      Out = In[OUT_SIZE*80-1:OUT_SIZE*79];
        7'd80:      Out = In[OUT_SIZE*81-1:OUT_SIZE*80];
        7'd81:      Out = In[OUT_SIZE*82-1:OUT_SIZE*81];
        7'd82:      Out = In[OUT_SIZE*83-1:OUT_SIZE*82];
        7'd83:      Out = In[OUT_SIZE*84-1:OUT_SIZE*83];
        7'd84:      Out = In[OUT_SIZE*85-1:OUT_SIZE*84];
        7'd85:      Out = In[OUT_SIZE*86-1:OUT_SIZE*85];
        7'd86:      Out = In[OUT_SIZE*87-1:OUT_SIZE*86];
        7'd87:      Out = In[OUT_SIZE*88-1:OUT_SIZE*87];
        7'd88:      Out = In[OUT_SIZE*89-1:OUT_SIZE*88];
        7'd89:      Out = In[OUT_SIZE*90-1:OUT_SIZE*89];
        7'd90:      Out = In[OUT_SIZE*91-1:OUT_SIZE*90];
        7'd91:      Out = In[OUT_SIZE*92-1:OUT_SIZE*91];
        7'd92:      Out = In[OUT_SIZE*93-1:OUT_SIZE*92];
        7'd93:      Out = In[OUT_SIZE*94-1:OUT_SIZE*93];
        7'd94:      Out = In[OUT_SIZE*95-1:OUT_SIZE*94];
        7'd95:      Out = In[OUT_SIZE*96-1:OUT_SIZE*95];
        7'd96:      Out = In[OUT_SIZE*97-1:OUT_SIZE*96];
        7'd97:      Out = In[OUT_SIZE*98-1:OUT_SIZE*97];
        7'd98:      Out = In[OUT_SIZE*99-1:OUT_SIZE*98];
        7'd99:      Out = In[OUT_SIZE*100-1:OUT_SIZE*99];
        7'd100:      Out = In[OUT_SIZE*101-1:OUT_SIZE*100];
        7'd101:      Out = In[OUT_SIZE*102-1:OUT_SIZE*101];
        7'd102:      Out = In[OUT_SIZE*103-1:OUT_SIZE*102];
        7'd103:      Out = In[OUT_SIZE*104-1:OUT_SIZE*103];
        7'd104:      Out = In[OUT_SIZE*105-1:OUT_SIZE*104];
        7'd105:      Out = In[OUT_SIZE*106-1:OUT_SIZE*105];
        7'd106:      Out = In[OUT_SIZE*107-1:OUT_SIZE*106];
        7'd107:      Out = In[OUT_SIZE*108-1:OUT_SIZE*107];
        7'd108:      Out = In[OUT_SIZE*109-1:OUT_SIZE*108];
        7'd109:      Out = In[OUT_SIZE*110-1:OUT_SIZE*109];
        7'd110:      Out = In[OUT_SIZE*111-1:OUT_SIZE*110];
        7'd111:      Out = In[OUT_SIZE*112-1:OUT_SIZE*111];
    endcase
end

endmodule
