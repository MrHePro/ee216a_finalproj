//TESTED
module Mux_Pixel(In, Select, Out);

parameter OUT_SIZE = 280;
parameter SEL_SIZE = 28;
parameter SEL_BIT  = 5;

input       [OUT_SIZE*SEL_SIZE-1:0]     In;
input       [SEL_BIT-1:0]               Select;
output  reg [OUT_SIZE-1:0]              Out;

always@(Select) begin
    case(Select)
        default:    Out = In[OUT_SIZE*1-1:OUT_SIZE*0];
        5'd1:       Out = In[OUT_SIZE*2-1:OUT_SIZE*1];
        5'd2:       Out = In[OUT_SIZE*3-1:OUT_SIZE*2];
        5'd3:       Out = In[OUT_SIZE*4-1:OUT_SIZE*3];
        5'd4:       Out = In[OUT_SIZE*5-1:OUT_SIZE*4];
        5'd5:       Out = In[OUT_SIZE*6-1:OUT_SIZE*5];
        5'd6:       Out = In[OUT_SIZE*7-1:OUT_SIZE*6];
        5'd7:       Out = In[OUT_SIZE*8-1:OUT_SIZE*7];
        5'd8:       Out = In[OUT_SIZE*9-1:OUT_SIZE*8];
        5'd9:       Out = In[OUT_SIZE*10-1:OUT_SIZE*9];
        5'd10:      Out = In[OUT_SIZE*11-1:OUT_SIZE*10];
        5'd11:      Out = In[OUT_SIZE*12-1:OUT_SIZE*11];
        5'd12:      Out = In[OUT_SIZE*13-1:OUT_SIZE*12];
        5'd13:      Out = In[OUT_SIZE*14-1:OUT_SIZE*13];
        5'd14:      Out = In[OUT_SIZE*15-1:OUT_SIZE*14];
        5'd15:      Out = In[OUT_SIZE*16-1:OUT_SIZE*15];
        5'd16:      Out = In[OUT_SIZE*17-1:OUT_SIZE*16];
        5'd17:      Out = In[OUT_SIZE*18-1:OUT_SIZE*17];
        5'd18:      Out = In[OUT_SIZE*19-1:OUT_SIZE*18];
        5'd19:      Out = In[OUT_SIZE*20-1:OUT_SIZE*19];
        5'd20:      Out = In[OUT_SIZE*21-1:OUT_SIZE*20];
        5'd21:      Out = In[OUT_SIZE*22-1:OUT_SIZE*21];
        5'd22:      Out = In[OUT_SIZE*23-1:OUT_SIZE*22];
        5'd23:      Out = In[OUT_SIZE*24-1:OUT_SIZE*23];
        5'd24:      Out = In[OUT_SIZE*25-1:OUT_SIZE*24];
        5'd25:      Out = In[OUT_SIZE*26-1:OUT_SIZE*25];
        5'd26:      Out = In[OUT_SIZE*27-1:OUT_SIZE*26];
        5'd27:      Out = In[OUT_SIZE*28-1:OUT_SIZE*27];
        5'd28:      Out = In[OUT_SIZE*29-1:OUT_SIZE*28];
        5'd29:      Out = In[OUT_SIZE*30-1:OUT_SIZE*29];
        5'd30:      Out = In[OUT_SIZE*31-1:OUT_SIZE*30];
        5'd31:      Out = In[OUT_SIZE*32-1:OUT_SIZE*31];
        5'd32:      Out = In[OUT_SIZE*33-1:OUT_SIZE*32];
        5'd33:      Out = In[OUT_SIZE*34-1:OUT_SIZE*33];
        5'd34:      Out = In[OUT_SIZE*35-1:OUT_SIZE*34];
        5'd35:      Out = In[OUT_SIZE*36-1:OUT_SIZE*35];
        5'd36:      Out = In[OUT_SIZE*37-1:OUT_SIZE*36];
        5'd37:      Out = In[OUT_SIZE*38-1:OUT_SIZE*37];
        5'd38:      Out = In[OUT_SIZE*39-1:OUT_SIZE*38];
        5'd39:      Out = In[OUT_SIZE*40-1:OUT_SIZE*39];
        5'd40:      Out = In[OUT_SIZE*41-1:OUT_SIZE*40];
        5'd41:      Out = In[OUT_SIZE*42-1:OUT_SIZE*41];
        5'd42:      Out = In[OUT_SIZE*43-1:OUT_SIZE*42];
        5'd43:      Out = In[OUT_SIZE*44-1:OUT_SIZE*43];
        5'd44:      Out = In[OUT_SIZE*45-1:OUT_SIZE*44];
        5'd45:      Out = In[OUT_SIZE*46-1:OUT_SIZE*45];
        5'd46:      Out = In[OUT_SIZE*47-1:OUT_SIZE*46];
        5'd47:      Out = In[OUT_SIZE*48-1:OUT_SIZE*47];
        5'd48:      Out = In[OUT_SIZE*49-1:OUT_SIZE*48];
        5'd49:      Out = In[OUT_SIZE*50-1:OUT_SIZE*49];
        5'd50:      Out = In[OUT_SIZE*51-1:OUT_SIZE*50];
        5'd51:      Out = In[OUT_SIZE*52-1:OUT_SIZE*51];
        5'd52:      Out = In[OUT_SIZE*53-1:OUT_SIZE*52];
        5'd53:      Out = In[OUT_SIZE*54-1:OUT_SIZE*53];
        5'd54:      Out = In[OUT_SIZE*55-1:OUT_SIZE*54];
        5'd55:      Out = In[OUT_SIZE*56-1:OUT_SIZE*55];
        5'd56:      Out = In[OUT_SIZE*57-1:OUT_SIZE*56];
        5'd57:      Out = In[OUT_SIZE*58-1:OUT_SIZE*57];
        5'd58:      Out = In[OUT_SIZE*59-1:OUT_SIZE*58];
        5'd59:      Out = In[OUT_SIZE*60-1:OUT_SIZE*59];
        5'd60:      Out = In[OUT_SIZE*61-1:OUT_SIZE*60];
        5'd61:      Out = In[OUT_SIZE*62-1:OUT_SIZE*61];
        5'd62:      Out = In[OUT_SIZE*63-1:OUT_SIZE*62];
        5'd63:      Out = In[OUT_SIZE*64-1:OUT_SIZE*63];
        5'd64:      Out = In[OUT_SIZE*65-1:OUT_SIZE*64];
        5'd65:      Out = In[OUT_SIZE*66-1:OUT_SIZE*65];
        5'd66:      Out = In[OUT_SIZE*67-1:OUT_SIZE*66];
        5'd67:      Out = In[OUT_SIZE*68-1:OUT_SIZE*67];
        5'd68:      Out = In[OUT_SIZE*69-1:OUT_SIZE*68];
        5'd69:      Out = In[OUT_SIZE*70-1:OUT_SIZE*69];
        5'd70:      Out = In[OUT_SIZE*71-1:OUT_SIZE*70];
        5'd71:      Out = In[OUT_SIZE*72-1:OUT_SIZE*71];
        5'd72:      Out = In[OUT_SIZE*73-1:OUT_SIZE*72];
        5'd73:      Out = In[OUT_SIZE*74-1:OUT_SIZE*73];
        5'd74:      Out = In[OUT_SIZE*75-1:OUT_SIZE*74];
        5'd75:      Out = In[OUT_SIZE*76-1:OUT_SIZE*75];
        5'd76:      Out = In[OUT_SIZE*77-1:OUT_SIZE*76];
        5'd77:      Out = In[OUT_SIZE*78-1:OUT_SIZE*77];
        5'd78:      Out = In[OUT_SIZE*79-1:OUT_SIZE*78];
        5'd79:      Out = In[OUT_SIZE*80-1:OUT_SIZE*79];
        5'd80:      Out = In[OUT_SIZE*81-1:OUT_SIZE*80];
        5'd81:      Out = In[OUT_SIZE*82-1:OUT_SIZE*81];
        5'd82:      Out = In[OUT_SIZE*83-1:OUT_SIZE*82];
        5'd83:      Out = In[OUT_SIZE*84-1:OUT_SIZE*83];
        5'd84:      Out = In[OUT_SIZE*85-1:OUT_SIZE*84];
        5'd85:      Out = In[OUT_SIZE*86-1:OUT_SIZE*85];
        5'd86:      Out = In[OUT_SIZE*87-1:OUT_SIZE*86];
        5'd87:      Out = In[OUT_SIZE*88-1:OUT_SIZE*87];
        5'd88:      Out = In[OUT_SIZE*89-1:OUT_SIZE*88];
        5'd89:      Out = In[OUT_SIZE*90-1:OUT_SIZE*89];
        5'd90:      Out = In[OUT_SIZE*91-1:OUT_SIZE*90];
        5'd91:      Out = In[OUT_SIZE*92-1:OUT_SIZE*91];
        5'd92:      Out = In[OUT_SIZE*93-1:OUT_SIZE*92];
        5'd93:      Out = In[OUT_SIZE*94-1:OUT_SIZE*93];
        5'd94:      Out = In[OUT_SIZE*95-1:OUT_SIZE*94];
        5'd95:      Out = In[OUT_SIZE*96-1:OUT_SIZE*95];
        5'd96:      Out = In[OUT_SIZE*97-1:OUT_SIZE*96];
        5'd97:      Out = In[OUT_SIZE*98-1:OUT_SIZE*97];
        5'd98:      Out = In[OUT_SIZE*99-1:OUT_SIZE*98];
        5'd99:      Out = In[OUT_SIZE*100-1:OUT_SIZE*99];
        5'd100:      Out = In[OUT_SIZE*101-1:OUT_SIZE*100];
        5'd101:      Out = In[OUT_SIZE*102-1:OUT_SIZE*101];
        5'd102:      Out = In[OUT_SIZE*103-1:OUT_SIZE*102];
        5'd103:      Out = In[OUT_SIZE*104-1:OUT_SIZE*103];
        5'd104:      Out = In[OUT_SIZE*105-1:OUT_SIZE*104];
        5'd105:      Out = In[OUT_SIZE*106-1:OUT_SIZE*105];
        5'd106:      Out = In[OUT_SIZE*107-1:OUT_SIZE*106];
        5'd107:      Out = In[OUT_SIZE*108-1:OUT_SIZE*107];
        5'd108:      Out = In[OUT_SIZE*109-1:OUT_SIZE*108];
        5'd109:      Out = In[OUT_SIZE*110-1:OUT_SIZE*109];
        5'd110:      Out = In[OUT_SIZE*111-1:OUT_SIZE*110];
        5'd111:      Out = In[OUT_SIZE*112-1:OUT_SIZE*111];
        5'd112:      Out = In[OUT_SIZE*113-1:OUT_SIZE*112];
    endcase
end

endmodule
